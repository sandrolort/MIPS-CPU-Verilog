module ff1_tb;
    parameter N = 32;
    reg [N-1:0] x;
    wire [4:0] y;

    ff1 #(N) uut (.x(x), .y(y));

    initial begin
        $monitor($time, " x = %b, y = %b", x, y);
        x = 32'b00000000000000000000000000000000; #10;
        x = 32'b10000000000000000000000000000000; #10;
        x = 32'b11000000000000000000000000000000; #10;
        x = 32'b11100000000000000000000000000000; #10;
        x = 32'b11111111000000000000000000000000; #10;
        x = 32'b10101010101010101010101010101010; #10;
        x = 32'b01010101010101010101010101010101; #10;
        x = 32'b00000000000000100000000000000000; #10;
        x = 32'b00000000100000000000000000000000; #10;
        x = 32'b00000000000000000010000000000000; #10;
        x = 32'b00000000000000000010000000000001; #10;
    end
endmodule
